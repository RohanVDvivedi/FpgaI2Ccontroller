
// The given main module, queries accelerometer data and gyroscope data, over i2c and 
module main(
    );


endmodule
